module d_fif_tb ;
    
    reg d,clk,rst;

    wire q;

    d_fif dut(
        .d(d),
        .clk(clk),
        .rst(rst),
        .q(q)
    );

    always #5 clk =~ clk;

    initial begin
        clk = 0;
        rst = 1;
        #5
        rst = 0;

        d = 0;
        #10 d = 1;
        #10 d = 0;
        #10 d = 1;
        #10 d = 0;
        #10 $finish;
    end

    initial begin
        $dumpfile("d_fif.vcd");
        $dumpvars(0,d_fif_tb);
    end
endmodule